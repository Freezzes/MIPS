library verilog;
use verilog.vl_types.all;
entity rtype_vlg_vec_tst is
end rtype_vlg_vec_tst;
